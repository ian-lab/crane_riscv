module rom (
    input [31:0] addr,
    output reg [31:0] instr
);

reg [31:0] rom [31:0];

// initial $readmemb("", bin_mem);
initial begin
  // Load instructions into ROM
  rom[0] = 32'b00000000000100000000000010010011; // addi x1, x0, 1
  rom[1] = 32'b00000000001000000000000100010011; // addi x2, x0, 2
  rom[2] = 32'b00000000001100000000000110010011; // addi x3, x0, 3
  rom[3] = 32'b00000000010000000000001000010011; // addi x4, x0, 4
  rom[4] = 32'b00000000010100000000001010010011; // addi x5, x0, 5
  rom[5] = 32'b00000000011000000000001100010011; // addi x6, x0, 6
  rom[6] = 32'b00000000011100000000001110010011; // addi x7, x0, 7
  rom[7] = 32'b00000000100000000000010000010011; // addi x8, x0, 8
  rom[8] = 32'b00000000100100000000010010010011; // addi x9, x0, 9
  rom[9] = 32'b00000000101000000000010100010011; // addi x10, x0, 10
  rom[10] = 32'b00000000101100000000010110010011; // addi x11, x0, 11
  rom[11] = 32'b00000000110000000000011000010011; // addi x12, x0, 12
end

always @(*) begin
    instr = rom[addr[31:2]];
    $display("rom[%d] = %h", addr[31:2], instr);
end
    
endmodule