module rom (
    input [31:0] addr,
    output reg [31:0] instr
);

reg [31:0] rom [31:0];

// initial $readmemb("", bin_mem);
initial begin
  rom[0] = 32'b0000_0000_0010_0001_0000_0010_1011_0011; // addi x2, x0, 2 hex: 0X002102B3
  rom[1] = 32'b0000_0000_0011_0001_0000_0011_1011_0011; // addi x3, x0, 3 hex: 0x003102B3
  rom[2] = 32'b0000_0000_0100_0001_0000_0100_1011_0011; // addi x4, x0, 4 hex: 0x004102B3
  rom[3] = 32'b0000_0000_0101_0001_0000_0101_1011_0011; // addi x5, x0, 5 hex: 0x005102B3
  rom[4] = 32'b0000_0000_0010_0001_0000_0010_1011_0011; // addi x2, x0, 2 
  rom[5] = 32'b0000_0000_0011_0001_0000_0011_1011_0011; // addi x3, x0, 3 
  rom[6] = 32'b0000_0000_0100_0001_0000_0100_1011_0011; // addi x4, x0, 4 
  rom[7] = 32'b0000_0000_0101_0001_0000_0101_1011_0011; // addi x5, x0, 5 
end

always @(*) begin
    instr = rom[addr[31:2]];
    $display("rom[%d] = %h", addr[31:2], instr);
end
    
endmodule